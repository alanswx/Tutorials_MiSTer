typedef enum bit[4:0] { 
BANK00, BANKF8, BANKF6, BANKFE, BANKE0, BANK3F, BANKF4, BANKP2, 
BANKFA, BANKCV, BANK2K, BANKUA, BANKE7, BANKF0, BANK32, BANKAR,
BANK3E, BANKSB, BANKWD, BANKEF, BANKDPCP, BANKCTY, BANKCDF
} bss_type ;

